VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AAOAOI33111
  CLASS CORE ;
  FOREIGN AAOAOI33111 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.300 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 12.300 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 12.300 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 11.650 3.150 12.150 3.650 ;
        RECT 11.750 2.300 12.050 3.150 ;
        RECT 11.650 1.800 12.150 2.300 ;
    END
  END Y
  PIN B2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 7.600 2.350 8.050 3.200 ;
    END
  END B2
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 9.850 2.350 10.300 3.200 ;
    END
  END A1
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 10.950 2.350 11.450 3.200 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.750 3.600 2.800 ;
        RECT 4.250 2.750 4.700 3.200 ;
        RECT 3.150 2.450 4.600 2.750 ;
        RECT 3.150 2.350 3.600 2.450 ;
    END
  END C
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.350 9.200 3.200 ;
    END
  END A2
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.350 2.350 5.850 3.200 ;
    END
  END B
  PIN B1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.500 2.350 6.950 3.200 ;
    END
  END B1
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.350 1.350 3.200 ;
    END
  END E
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 1.750 2.350 2.200 2.800 ;
    END
  END D
END AAOAOI33111
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND4
  CLASS CORE ;
  FOREIGN NAND4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.600 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 5.600 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 5.600 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.200 3.550 0.650 3.650 ;
        RECT 4.950 3.550 5.400 3.650 ;
        RECT 0.200 3.250 5.400 3.550 ;
        RECT 0.200 3.150 0.650 3.250 ;
        RECT 4.950 3.150 5.400 3.250 ;
        RECT 5.050 2.300 5.300 3.150 ;
        RECT 4.950 1.800 5.400 2.300 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.250 2.350 4.700 2.800 ;
    END
  END A
  PIN A3
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.350 1.350 2.800 ;
    END
  END A3
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.350 3.600 2.800 ;
    END
  END A1
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 2.350 2.450 2.800 ;
    END
  END A2
END NAND4
END LIBRARY


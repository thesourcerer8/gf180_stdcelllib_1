VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO AAAOAI3221
  CLASS CORE ;
  FOREIGN AAAOAI3221 ;
  ORIGIN 0.000 0.000 ;
  SIZE 11.200 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 11.200 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 11.200 0.250 ;
    END
  END VGND
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 10.550 3.150 11.000 3.650 ;
        RECT 10.650 2.300 10.900 3.150 ;
        RECT 10.550 1.800 11.000 2.300 ;
    END
  END Y
  PIN A2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 7.600 2.350 8.050 3.200 ;
    END
  END A2
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 9.850 2.350 10.300 3.200 ;
    END
  END A
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.350 3.600 3.200 ;
    END
  END C
  PIN B1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.500 2.350 6.950 3.200 ;
    END
  END B1
  PIN A1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.350 9.200 3.200 ;
    END
  END A1
  PIN C1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 2.350 2.450 3.200 ;
    END
  END C1
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.350 2.350 5.850 3.200 ;
    END
  END B
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.350 1.350 3.200 ;
    END
  END D
END AAAOAI3221
END LIBRARY


MACRO AOAAOI2124
 CLASS CORE ;
 FOREIGN AOAAOI2124 0 0 ;
 SIZE 12.32 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 12.32000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 12.32000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 11.53000000 0.46700000 11.99000000 0.92700000 ;
    END
  END Y

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
    END
  END C1

  PIN D1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
    END
  END D1

  PIN D2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
    END
  END D2

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
    END
  END D

  PIN D3
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
    END
  END D3

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.10000000 2.17700000 11.34000000 2.35700000 ;
        RECT 9.10000000 2.35700000 11.43000000 2.45700000 ;
        RECT 9.10000000 2.45700000 9.38000000 2.76200000 ;
        RECT 10.97000000 2.45700000 11.43000000 2.81700000 ;
        RECT 9.01000000 2.76200000 9.47000000 3.22200000 ;
    END
  END A

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.85000000 2.76200000 10.31000000 3.22200000 ;
    END
  END A1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
    END
  END B

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 7.73000000 2.47700000 7.95000000 2.69700000 ;
     RECT 9.97000000 2.47700000 10.19000000 2.69700000 ;
     RECT 11.09000000 2.47700000 11.31000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;
     RECT 8.85000000 2.88200000 9.07000000 3.10200000 ;
     RECT 9.97000000 2.88200000 10.19000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.29500000 3.27200000 0.54500000 3.52200000 ;
     RECT 10.65500000 3.54200000 10.90500000 3.79200000 ;

    LAYER ndiffc ;
     RECT 4.91500000 0.30200000 5.16500000 0.55200000 ;
     RECT 7.15500000 0.57200000 7.40500000 0.82200000 ;
     RECT 9.25500000 0.57200000 9.50500000 0.82200000 ;
     RECT 11.63500000 0.57200000 11.88500000 0.82200000 ;
     RECT 0.29500000 1.92200000 0.54500000 2.17200000 ;
     RECT 8.41500000 1.92200000 8.66500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 12.32000000 0.24000000 ;
     RECT 4.83500000 0.24000000 5.24500000 0.63200000 ;
     RECT 7.07500000 0.49200000 7.48500000 0.90200000 ;
     RECT 9.17500000 0.49200000 9.58500000 0.90200000 ;
     RECT 11.55500000 0.49200000 11.96500000 0.90200000 ;
     RECT 0.21500000 1.84200000 0.62500000 2.25200000 ;
     RECT 8.33500000 1.84200000 8.74500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 4.29000000 2.39700000 4.67000000 2.77700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 7.65000000 2.39700000 8.03000000 2.77700000 ;
     RECT 11.01000000 2.39700000 11.39000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.80200000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.80200000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.80200000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.80200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.80200000 9.43000000 3.18200000 ;
     RECT 9.89000000 2.39700000 10.27000000 3.18200000 ;
     RECT 0.21500000 3.19200000 0.62500000 3.60200000 ;
     RECT 10.57500000 3.46200000 10.98500000 3.87200000 ;
     RECT 0.00000000 4.80000000 12.32000000 5.28000000 ;

    LAYER via1 ;
     RECT 7.15000000 0.56700000 7.41000000 0.82700000 ;
     RECT 9.25000000 0.56700000 9.51000000 0.82700000 ;
     RECT 11.63000000 0.56700000 11.89000000 0.82700000 ;
     RECT 0.29000000 1.91700000 0.55000000 2.17700000 ;
     RECT 8.41000000 1.91700000 8.67000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 4.35000000 2.45700000 4.61000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 7.71000000 2.45700000 7.97000000 2.71700000 ;
     RECT 11.07000000 2.45700000 11.33000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 2.86200000 2.37000000 3.12200000 ;
     RECT 3.23000000 2.86200000 3.49000000 3.12200000 ;
     RECT 4.35000000 2.86200000 4.61000000 3.12200000 ;
     RECT 5.47000000 2.86200000 5.73000000 3.12200000 ;
     RECT 6.59000000 2.86200000 6.85000000 3.12200000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 9.11000000 2.86200000 9.37000000 3.12200000 ;
     RECT 9.95000000 2.86200000 10.21000000 3.12200000 ;
     RECT 0.29000000 3.26700000 0.55000000 3.52700000 ;
     RECT 10.65000000 3.53700000 10.91000000 3.79700000 ;

    LAYER met2 ;
     RECT 7.05000000 0.46700000 7.51000000 0.55700000 ;
     RECT 9.15000000 0.46700000 9.61000000 0.55700000 ;
     RECT 7.05000000 0.55700000 9.61000000 0.83700000 ;
     RECT 7.05000000 0.83700000 7.51000000 0.92700000 ;
     RECT 9.15000000 0.83700000 9.61000000 0.92700000 ;
     RECT 11.53000000 0.46700000 11.99000000 0.92700000 ;
     RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
     RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
     RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
     RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
     RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
     RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
     RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
     RECT 9.10000000 2.17700000 11.34000000 2.35700000 ;
     RECT 9.10000000 2.35700000 11.43000000 2.45700000 ;
     RECT 9.10000000 2.45700000 9.38000000 2.76200000 ;
     RECT 10.97000000 2.45700000 11.43000000 2.81700000 ;
     RECT 9.01000000 2.76200000 9.47000000 3.22200000 ;
     RECT 9.85000000 2.76200000 10.31000000 3.22200000 ;
     RECT 0.19000000 1.81700000 0.65000000 2.27700000 ;
     RECT 0.28000000 2.27700000 0.56000000 3.16700000 ;
     RECT 0.19000000 3.16700000 0.65000000 3.62700000 ;
     RECT 8.31000000 1.81700000 8.77000000 2.27700000 ;
     RECT 8.40000000 2.27700000 8.68000000 3.52700000 ;
     RECT 10.55000000 3.43700000 11.01000000 3.52700000 ;
     RECT 8.40000000 3.52700000 11.01000000 3.80700000 ;
     RECT 10.55000000 3.80700000 11.01000000 3.89700000 ;

 END
END AOAAOI2124

MACRO ASYNC3
 CLASS CORE ;
 FOREIGN ASYNC3 0 0 ;
 SIZE 8.96 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 8.96000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 8.96000000 0.24000000 ;
    END
  END GND

  PIN CN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 1.45000000 1.68200000 1.91000000 1.77200000 ;
        RECT 7.61000000 1.68200000 8.07000000 1.77200000 ;
        RECT 1.45000000 1.77200000 8.07000000 2.05200000 ;
        RECT 1.45000000 2.05200000 1.91000000 2.14200000 ;
        RECT 7.61000000 2.05200000 8.07000000 2.14200000 ;
    END
  END CN

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 8.31000000 1.81700000 8.77000000 2.27700000 ;
        RECT 5.37000000 2.35700000 5.83000000 2.44700000 ;
        RECT 8.40000000 2.27700000 8.68000000 2.44700000 ;
        RECT 5.37000000 2.44700000 8.68000000 2.72700000 ;
        RECT 5.37000000 2.72700000 5.83000000 2.81700000 ;
        RECT 8.40000000 2.72700000 8.68000000 3.16700000 ;
        RECT 8.31000000 3.16700000 8.77000000 3.62700000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 2.44700000 ;
        RECT 3.13000000 2.35700000 3.59000000 2.44700000 ;
        RECT 0.89000000 2.44700000 3.59000000 2.72700000 ;
        RECT 3.13000000 2.72700000 3.59000000 2.81700000 ;
        RECT 0.89000000 2.72700000 1.35000000 3.22200000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.01000000 3.03200000 2.47000000 3.12200000 ;
        RECT 6.49000000 3.03200000 6.95000000 3.12200000 ;
        RECT 2.01000000 3.12200000 6.95000000 3.40200000 ;
        RECT 2.01000000 3.40200000 2.47000000 3.49200000 ;
        RECT 6.49000000 3.40200000 6.95000000 3.49200000 ;
    END
  END B

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 7.73000000 2.47700000 7.95000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 8.41500000 3.27200000 8.66500000 3.52200000 ;
     RECT 3.93500000 4.48700000 4.18500000 4.73700000 ;

    LAYER ndiffc ;
     RECT 3.79500000 0.30200000 4.04500000 0.55200000 ;
     RECT 7.15500000 0.30200000 7.40500000 0.55200000 ;
     RECT 0.43500000 0.57200000 0.68500000 0.82200000 ;
     RECT 6.03500000 0.57200000 6.28500000 0.82200000 ;
     RECT 2.67500000 0.70700000 2.92500000 0.95700000 ;
     RECT 4.77500000 0.70700000 5.02500000 0.95700000 ;
     RECT 1.55500000 1.78700000 1.80500000 2.03700000 ;
     RECT 8.41500000 1.92200000 8.66500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 8.96000000 0.24000000 ;
     RECT 3.71500000 0.24000000 4.12500000 0.63200000 ;
     RECT 7.07500000 0.24000000 7.48500000 0.63200000 ;
     RECT 0.35500000 0.49200000 0.76500000 0.90200000 ;
     RECT 5.95500000 0.49200000 6.36500000 0.90200000 ;
     RECT 2.59500000 0.62700000 3.00500000 1.03700000 ;
     RECT 4.69500000 0.62700000 5.10500000 1.03700000 ;
     RECT 1.47500000 1.70700000 1.88500000 2.11700000 ;
     RECT 8.33500000 1.84200000 8.74500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;
     RECT 5.41000000 2.39700000 5.79000000 3.18200000 ;
     RECT 7.65000000 1.72200000 8.03000000 2.10200000 ;
     RECT 7.72500000 2.10200000 7.95500000 2.39700000 ;
     RECT 7.65000000 2.39700000 8.03000000 3.18200000 ;
     RECT 2.05000000 2.39700000 2.43000000 3.45200000 ;
     RECT 6.53000000 2.39700000 6.91000000 3.45200000 ;
     RECT 8.33500000 3.19200000 8.74500000 3.60200000 ;
     RECT 3.85500000 4.40700000 4.26500000 4.80000000 ;
     RECT 0.00000000 4.80000000 8.96000000 5.28000000 ;

    LAYER via1 ;
     RECT 0.43000000 0.56700000 0.69000000 0.82700000 ;
     RECT 6.03000000 0.56700000 6.29000000 0.82700000 ;
     RECT 2.67000000 0.70200000 2.93000000 0.96200000 ;
     RECT 4.77000000 0.70200000 5.03000000 0.96200000 ;
     RECT 1.55000000 1.78200000 1.81000000 2.04200000 ;
     RECT 7.71000000 1.78200000 7.97000000 2.04200000 ;
     RECT 8.41000000 1.91700000 8.67000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 3.13200000 2.37000000 3.39200000 ;
     RECT 6.59000000 3.13200000 6.85000000 3.39200000 ;
     RECT 8.41000000 3.26700000 8.67000000 3.52700000 ;

    LAYER met2 ;
     RECT 0.42000000 0.01700000 6.30000000 0.29700000 ;
     RECT 0.42000000 0.29700000 0.70000000 0.46700000 ;
     RECT 6.02000000 0.29700000 6.30000000 0.46700000 ;
     RECT 0.33000000 0.46700000 0.79000000 0.92700000 ;
     RECT 5.93000000 0.46700000 6.39000000 0.92700000 ;
     RECT 2.57000000 0.60200000 3.03000000 0.69200000 ;
     RECT 4.67000000 0.60200000 5.13000000 0.69200000 ;
     RECT 2.57000000 0.69200000 5.13000000 0.97200000 ;
     RECT 2.57000000 0.97200000 3.03000000 1.06200000 ;
     RECT 4.67000000 0.97200000 5.13000000 1.06200000 ;
     RECT 1.45000000 1.68200000 1.91000000 1.77200000 ;
     RECT 7.61000000 1.68200000 8.07000000 1.77200000 ;
     RECT 1.45000000 1.77200000 8.07000000 2.05200000 ;
     RECT 1.45000000 2.05200000 1.91000000 2.14200000 ;
     RECT 7.61000000 2.05200000 8.07000000 2.14200000 ;
     RECT 0.89000000 2.35700000 1.35000000 2.44700000 ;
     RECT 3.13000000 2.35700000 3.59000000 2.44700000 ;
     RECT 0.89000000 2.44700000 3.59000000 2.72700000 ;
     RECT 3.13000000 2.72700000 3.59000000 2.81700000 ;
     RECT 0.89000000 2.72700000 1.35000000 3.22200000 ;
     RECT 2.01000000 3.03200000 2.47000000 3.12200000 ;
     RECT 6.49000000 3.03200000 6.95000000 3.12200000 ;
     RECT 2.01000000 3.12200000 6.95000000 3.40200000 ;
     RECT 2.01000000 3.40200000 2.47000000 3.49200000 ;
     RECT 6.49000000 3.40200000 6.95000000 3.49200000 ;
     RECT 8.31000000 1.81700000 8.77000000 2.27700000 ;
     RECT 5.37000000 2.35700000 5.83000000 2.44700000 ;
     RECT 8.40000000 2.27700000 8.68000000 2.44700000 ;
     RECT 5.37000000 2.44700000 8.68000000 2.72700000 ;
     RECT 5.37000000 2.72700000 5.83000000 2.81700000 ;
     RECT 8.40000000 2.72700000 8.68000000 3.16700000 ;
     RECT 8.31000000 3.16700000 8.77000000 3.62700000 ;

 END
END ASYNC3

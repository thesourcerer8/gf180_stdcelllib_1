MACRO AAOAOI33111
 CLASS CORE ;
 FOREIGN AAOAOI33111 0 0 ;
 SIZE 12.32 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 12.32000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 12.32000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 11.67000000 1.81700000 12.13000000 2.27700000 ;
        RECT 11.76000000 2.27700000 12.04000000 3.16700000 ;
        RECT 11.67000000 3.16700000 12.13000000 3.62700000 ;
    END
  END Y

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
    END
  END B2

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.85000000 2.35700000 10.31000000 3.22200000 ;
    END
  END A1

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 10.97000000 2.35700000 11.43000000 3.22200000 ;
    END
  END A

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.13000000 2.35700000 3.59000000 2.44700000 ;
        RECT 3.13000000 2.44700000 4.62000000 2.72700000 ;
        RECT 4.25000000 2.72700000 4.62000000 2.76200000 ;
        RECT 3.13000000 2.72700000 3.59000000 2.81700000 ;
        RECT 4.25000000 2.76200000 4.71000000 3.22200000 ;
    END
  END C

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 8.73000000 2.35700000 9.19000000 3.22200000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
    END
  END B

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
    END
  END B1

  PIN E
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
    END
  END E

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 1.73000000 2.35700000 2.19000000 2.81700000 ;
    END
  END D

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 7.73000000 2.47700000 7.95000000 2.69700000 ;
     RECT 8.85000000 2.47700000 9.07000000 2.69700000 ;
     RECT 9.97000000 2.47700000 10.19000000 2.69700000 ;
     RECT 11.09000000 2.47700000 11.31000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;
     RECT 8.85000000 2.88200000 9.07000000 3.10200000 ;
     RECT 9.97000000 2.88200000 10.19000000 3.10200000 ;
     RECT 11.09000000 2.88200000 11.31000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 11.77500000 3.27200000 12.02500000 3.52200000 ;
     RECT 2.81500000 3.54200000 3.06500000 3.79200000 ;
     RECT 3.65500000 4.21700000 3.90500000 4.46700000 ;
     RECT 0.29500000 4.48700000 0.54500000 4.73700000 ;

    LAYER ndiffc ;
     RECT 1.55500000 0.30200000 1.80500000 0.55200000 ;
     RECT 2.67500000 0.57200000 2.92500000 0.82200000 ;
     RECT 8.27500000 0.57200000 8.52500000 0.82200000 ;
     RECT 0.29500000 1.92200000 0.54500000 2.17200000 ;
     RECT 11.77500000 1.92200000 12.02500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 12.32000000 0.24000000 ;
     RECT 1.47500000 0.24000000 1.88500000 0.63200000 ;
     RECT 2.59500000 0.49200000 3.00500000 0.90200000 ;
     RECT 8.19500000 0.49200000 8.60500000 0.90200000 ;
     RECT 0.21500000 1.84200000 0.62500000 2.25200000 ;
     RECT 11.69500000 1.84200000 12.10500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 7.65000000 2.39700000 8.03000000 2.77700000 ;
     RECT 8.77000000 2.39700000 9.15000000 2.77700000 ;
     RECT 9.89000000 2.39700000 10.27000000 2.77700000 ;
     RECT 11.01000000 2.39700000 11.39000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 1.77000000 2.39700000 2.43000000 2.77700000 ;
     RECT 2.05000000 2.77700000 2.43000000 3.18200000 ;
     RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.80200000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.80200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.80200000 9.15000000 3.18200000 ;
     RECT 9.89000000 2.80200000 10.27000000 3.18200000 ;
     RECT 11.01000000 2.80200000 11.39000000 3.18200000 ;
     RECT 11.69500000 3.19200000 12.10500000 3.60200000 ;
     RECT 2.73500000 3.46200000 3.14500000 3.87200000 ;
     RECT 3.57500000 4.13700000 3.98500000 4.54700000 ;
     RECT 0.21500000 4.40700000 0.62500000 4.80000000 ;
     RECT 0.00000000 4.80000000 12.32000000 5.28000000 ;

    LAYER via1 ;
     RECT 2.67000000 0.56700000 2.93000000 0.82700000 ;
     RECT 8.27000000 0.56700000 8.53000000 0.82700000 ;
     RECT 0.29000000 1.91700000 0.55000000 2.17700000 ;
     RECT 11.77000000 1.91700000 12.03000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 1.83000000 2.45700000 2.09000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 7.71000000 2.45700000 7.97000000 2.71700000 ;
     RECT 8.83000000 2.45700000 9.09000000 2.71700000 ;
     RECT 9.95000000 2.45700000 10.21000000 2.71700000 ;
     RECT 11.07000000 2.45700000 11.33000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 4.35000000 2.86200000 4.61000000 3.12200000 ;
     RECT 5.47000000 2.86200000 5.73000000 3.12200000 ;
     RECT 6.59000000 2.86200000 6.85000000 3.12200000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 8.83000000 2.86200000 9.09000000 3.12200000 ;
     RECT 9.95000000 2.86200000 10.21000000 3.12200000 ;
     RECT 11.07000000 2.86200000 11.33000000 3.12200000 ;
     RECT 11.77000000 3.26700000 12.03000000 3.52700000 ;
     RECT 2.81000000 3.53700000 3.07000000 3.79700000 ;
     RECT 3.65000000 4.21200000 3.91000000 4.47200000 ;

    LAYER met2 ;
     RECT 1.73000000 2.35700000 2.19000000 2.81700000 ;
     RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
     RECT 3.13000000 2.35700000 3.59000000 2.44700000 ;
     RECT 3.13000000 2.44700000 4.62000000 2.72700000 ;
     RECT 4.25000000 2.72700000 4.62000000 2.76200000 ;
     RECT 3.13000000 2.72700000 3.59000000 2.81700000 ;
     RECT 4.25000000 2.76200000 4.71000000 3.22200000 ;
     RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
     RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
     RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
     RECT 8.73000000 2.35700000 9.19000000 3.22200000 ;
     RECT 9.85000000 2.35700000 10.31000000 3.22200000 ;
     RECT 10.97000000 2.35700000 11.43000000 3.22200000 ;
     RECT 11.67000000 1.81700000 12.13000000 2.27700000 ;
     RECT 11.76000000 2.27700000 12.04000000 3.16700000 ;
     RECT 11.67000000 3.16700000 12.13000000 3.62700000 ;
     RECT 2.57000000 0.46700000 3.03000000 0.55700000 ;
     RECT 8.17000000 0.46700000 8.63000000 0.55700000 ;
     RECT 2.52000000 0.55700000 8.63000000 0.83700000 ;
     RECT 2.52000000 0.83700000 3.03000000 0.92700000 ;
     RECT 8.17000000 0.83700000 8.63000000 0.92700000 ;
     RECT 2.52000000 0.92700000 2.80000000 3.43700000 ;
     RECT 2.52000000 3.43700000 3.17000000 3.80700000 ;
     RECT 2.71000000 3.80700000 3.17000000 3.89700000 ;
     RECT 0.19000000 1.81700000 0.65000000 2.27700000 ;
     RECT 0.28000000 2.27700000 0.56000000 4.20200000 ;
     RECT 3.55000000 4.11200000 4.01000000 4.20200000 ;
     RECT 0.28000000 4.20200000 4.01000000 4.48200000 ;
     RECT 3.55000000 4.48200000 4.01000000 4.57200000 ;

 END
END AAOAOI33111

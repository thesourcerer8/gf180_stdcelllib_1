MACRO AAOI22
 CLASS CORE ;
 FOREIGN AAOI22 0 0 ;
 SIZE 5.6000000000000005 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 5.60000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 5.60000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.81000000 0.46700000 5.27000000 0.92700000 ;
    END
  END Y

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.13000000 2.35700000 3.59000000 2.81700000 ;
    END
  END A1

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.25000000 2.35700000 4.71000000 2.81700000 ;
    END
  END A

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.01000000 2.35700000 2.47000000 2.81700000 ;
    END
  END B1

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 2.81700000 ;
    END
  END B

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.29500000 3.27200000 0.54500000 3.52200000 ;
     RECT 5.05500000 3.27200000 5.30500000 3.52200000 ;

    LAYER ndiffc ;
     RECT 2.67500000 0.30200000 2.92500000 0.55200000 ;
     RECT 4.91500000 0.57200000 5.16500000 0.82200000 ;
     RECT 0.29500000 1.92200000 0.54500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 5.60000000 0.24000000 ;
     RECT 2.59500000 0.24000000 3.00500000 0.63200000 ;
     RECT 4.83500000 0.49200000 5.24500000 0.90200000 ;
     RECT 0.21500000 1.84200000 0.62500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.39700000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.39700000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.39700000 4.67000000 3.18200000 ;
     RECT 0.21500000 3.19200000 0.62500000 3.60200000 ;
     RECT 4.97500000 3.19200000 5.38500000 3.60200000 ;
     RECT 0.00000000 4.80000000 5.60000000 5.28000000 ;

    LAYER via1 ;
     RECT 4.91000000 0.56700000 5.17000000 0.82700000 ;
     RECT 0.29000000 1.91700000 0.55000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 4.35000000 2.45700000 4.61000000 2.71700000 ;
     RECT 0.29000000 3.26700000 0.55000000 3.52700000 ;
     RECT 5.05000000 3.26700000 5.31000000 3.52700000 ;

    LAYER met2 ;
     RECT 4.81000000 0.46700000 5.27000000 0.92700000 ;
     RECT 0.89000000 2.35700000 1.35000000 2.81700000 ;
     RECT 2.01000000 2.35700000 2.47000000 2.81700000 ;
     RECT 3.13000000 2.35700000 3.59000000 2.81700000 ;
     RECT 4.25000000 2.35700000 4.71000000 2.81700000 ;
     RECT 0.19000000 1.81700000 0.65000000 2.27700000 ;
     RECT 0.28000000 2.27700000 0.56000000 3.16700000 ;
     RECT 0.19000000 3.16700000 0.65000000 3.25700000 ;
     RECT 4.95000000 3.16700000 5.41000000 3.25700000 ;
     RECT 0.19000000 3.25700000 5.41000000 3.53700000 ;
     RECT 0.19000000 3.53700000 0.65000000 3.62700000 ;
     RECT 4.95000000 3.53700000 5.41000000 3.62700000 ;

 END
END AAOI22

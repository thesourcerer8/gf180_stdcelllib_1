MACRO AAAAOI3322
 CLASS CORE ;
 FOREIGN AAAAOI3322 0 0 ;
 SIZE 13.44 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 13.44000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 13.44000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.19000000 1.81700000 0.65000000 2.27700000 ;
        RECT 0.28000000 2.27700000 0.56000000 3.16700000 ;
        RECT 0.19000000 3.16700000 0.65000000 3.62700000 ;
    END
  END Y

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 8.73000000 3.03200000 9.19000000 3.49200000 ;
    END
  END D

  PIN C1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 10.97000000 3.03200000 11.43000000 3.49200000 ;
    END
  END C1

  PIN B2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
    END
  END B2

  PIN B1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
    END
  END B1

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 12.09000000 2.35700000 12.55000000 2.44700000 ;
        RECT 7.70000000 2.44700000 12.55000000 2.72700000 ;
        RECT 7.70000000 2.72700000 8.07000000 2.76200000 ;
        RECT 12.09000000 2.72700000 12.55000000 2.81700000 ;
        RECT 7.61000000 2.76200000 8.07000000 3.22200000 ;
    END
  END C

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
    END
  END A

  PIN A2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
    END
  END A2

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
    END
  END B

  PIN A1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
    END
  END A1

  PIN D1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.85000000 3.03200000 10.31000000 3.49200000 ;
    END
  END D1

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 8.85000000 2.47700000 9.07000000 2.69700000 ;
     RECT 9.97000000 2.47700000 10.19000000 2.69700000 ;
     RECT 11.09000000 2.47700000 11.31000000 2.69700000 ;
     RECT 12.21000000 2.47700000 12.43000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;
     RECT 8.85000000 2.88200000 9.07000000 3.10200000 ;
     RECT 9.97000000 2.88200000 10.19000000 3.10200000 ;
     RECT 11.09000000 2.88200000 11.31000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 0.29500000 3.27200000 0.54500000 3.52200000 ;
     RECT 11.77500000 3.27200000 12.02500000 3.52200000 ;

    LAYER ndiffc ;
     RECT 3.79500000 0.30200000 4.04500000 0.55200000 ;
     RECT 10.51500000 0.30200000 10.76500000 0.55200000 ;
     RECT 0.29500000 1.92200000 0.54500000 2.17200000 ;
     RECT 12.89500000 1.92200000 13.14500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 13.44000000 0.24000000 ;
     RECT 3.71500000 0.24000000 4.12500000 0.63200000 ;
     RECT 10.43500000 0.24000000 10.84500000 0.63200000 ;
     RECT 0.21500000 1.84200000 0.62500000 2.25200000 ;
     RECT 12.81500000 1.84200000 13.22500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 4.29000000 2.39700000 4.67000000 2.77700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 12.13000000 2.39700000 12.51000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.80200000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.80200000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.80200000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.80200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.39700000 9.15000000 3.45200000 ;
     RECT 9.89000000 2.39700000 10.27000000 3.45200000 ;
     RECT 11.01000000 2.39700000 11.39000000 3.45200000 ;
     RECT 0.21500000 3.19200000 0.62500000 3.60200000 ;
     RECT 11.69500000 3.19200000 12.10500000 3.60200000 ;
     RECT 0.00000000 4.80000000 13.44000000 5.28000000 ;

    LAYER via1 ;
     RECT 0.29000000 1.91700000 0.55000000 2.17700000 ;
     RECT 12.89000000 1.91700000 13.15000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 4.35000000 2.45700000 4.61000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 12.19000000 2.45700000 12.45000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 2.86200000 2.37000000 3.12200000 ;
     RECT 3.23000000 2.86200000 3.49000000 3.12200000 ;
     RECT 4.35000000 2.86200000 4.61000000 3.12200000 ;
     RECT 5.47000000 2.86200000 5.73000000 3.12200000 ;
     RECT 6.59000000 2.86200000 6.85000000 3.12200000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 8.83000000 3.13200000 9.09000000 3.39200000 ;
     RECT 9.95000000 3.13200000 10.21000000 3.39200000 ;
     RECT 11.07000000 3.13200000 11.33000000 3.39200000 ;
     RECT 0.29000000 3.26700000 0.55000000 3.52700000 ;
     RECT 11.77000000 3.26700000 12.03000000 3.52700000 ;

    LAYER met2 ;
     RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
     RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
     RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
     RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
     RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
     RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
     RECT 12.09000000 2.35700000 12.55000000 2.44700000 ;
     RECT 7.70000000 2.44700000 12.55000000 2.72700000 ;
     RECT 7.70000000 2.72700000 8.07000000 2.76200000 ;
     RECT 12.09000000 2.72700000 12.55000000 2.81700000 ;
     RECT 7.61000000 2.76200000 8.07000000 3.22200000 ;
     RECT 8.73000000 3.03200000 9.19000000 3.49200000 ;
     RECT 9.85000000 3.03200000 10.31000000 3.49200000 ;
     RECT 10.97000000 3.03200000 11.43000000 3.49200000 ;
     RECT 0.19000000 1.81700000 0.65000000 2.27700000 ;
     RECT 0.28000000 2.27700000 0.56000000 3.16700000 ;
     RECT 0.19000000 3.16700000 0.65000000 3.62700000 ;
     RECT 12.79000000 1.81700000 13.25000000 2.27700000 ;
     RECT 11.67000000 3.16700000 12.13000000 3.25700000 ;
     RECT 12.88000000 2.27700000 13.16000000 3.25700000 ;
     RECT 11.67000000 3.25700000 13.16000000 3.53700000 ;
     RECT 11.67000000 3.53700000 12.13000000 3.62700000 ;

 END
END AAAAOI3322

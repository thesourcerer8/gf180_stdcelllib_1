MACRO INV
 CLASS CORE ;
 FOREIGN INV 0 0 ;
 SIZE 2.24 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 2.24000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 2.24000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 1.59000000 1.81700000 2.05000000 2.27700000 ;
        RECT 1.68000000 2.27700000 1.96000000 3.16700000 ;
        RECT 1.59000000 3.16700000 2.05000000 3.62700000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
    END
  END A

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 1.69500000 3.27200000 1.94500000 3.52200000 ;
     RECT 0.29500000 4.48700000 0.54500000 4.73700000 ;

    LAYER ndiffc ;
     RECT 0.29500000 0.30200000 0.54500000 0.55200000 ;
     RECT 1.69500000 1.92200000 1.94500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 2.24000000 0.24000000 ;
     RECT 0.21500000 0.24000000 0.62500000 0.63200000 ;
     RECT 1.61500000 1.84200000 2.02500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 1.61500000 3.19200000 2.02500000 3.60200000 ;
     RECT 0.21500000 4.40700000 0.62500000 4.80000000 ;
     RECT 0.00000000 4.80000000 2.24000000 5.28000000 ;

    LAYER via1 ;
     RECT 1.69000000 1.91700000 1.95000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 1.69000000 3.26700000 1.95000000 3.52700000 ;

    LAYER met2 ;
     RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
     RECT 1.59000000 1.81700000 2.05000000 2.27700000 ;
     RECT 1.68000000 2.27700000 1.96000000 3.16700000 ;
     RECT 1.59000000 3.16700000 2.05000000 3.62700000 ;

 END
END INV

MACRO MUX8
 CLASS CORE ;
 FOREIGN MUX8 0 0 ;
 SIZE 20.16 BY 5.04 ;
 ORIGIN 0 0 ;
 SYMMETRY X Y R90 ;
 SITE unit ;
  PIN VDD
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 4.80000000 20.16000000 5.28000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE POWER ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met1 ;
        RECT 0.00000000 -0.24000000 20.16000000 0.24000000 ;
    END
  END GND

  PIN Z
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 19.51000000 1.81700000 19.97000000 2.27700000 ;
        RECT 19.60000000 2.27700000 19.88000000 3.16700000 ;
        RECT 19.51000000 3.16700000 19.97000000 3.62700000 ;
    END
  END Z

  PIN IN4
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 13.21000000 2.35700000 13.67000000 3.22200000 ;
    END
  END IN4

  PIN S0
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
    END
  END S0

  PIN IN0
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
    END
  END IN0

  PIN S5
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 15.45000000 2.35700000 15.91000000 3.22200000 ;
    END
  END S5

  PIN S7
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
    END
  END S7

  PIN IN5
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 14.33000000 2.35700000 14.79000000 3.22200000 ;
    END
  END IN5

  PIN IN1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 8.73000000 2.35700000 9.19000000 3.22200000 ;
    END
  END IN1

  PIN S1
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
    END
  END S1

  PIN S3
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
    END
  END S3

  PIN S6
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 10.97000000 2.35700000 11.43000000 3.22200000 ;
    END
  END S6

  PIN S2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 16.57000000 2.35700000 17.03000000 3.22200000 ;
    END
  END S2

  PIN IN2
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 17.69000000 2.35700000 18.15000000 3.22200000 ;
    END
  END IN2

  PIN IN3
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
    END
  END IN3

  PIN IN7
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
    END
  END IN7

  PIN S4
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 12.09000000 2.35700000 12.55000000 3.22200000 ;
    END
  END S4

  PIN IN6
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 9.85000000 2.35700000 10.31000000 3.22200000 ;
    END
  END IN6

 OBS
    LAYER polycont ;
     RECT 1.01000000 2.47700000 1.23000000 2.69700000 ;
     RECT 2.13000000 2.47700000 2.35000000 2.69700000 ;
     RECT 3.25000000 2.47700000 3.47000000 2.69700000 ;
     RECT 4.37000000 2.47700000 4.59000000 2.69700000 ;
     RECT 5.49000000 2.47700000 5.71000000 2.69700000 ;
     RECT 6.61000000 2.47700000 6.83000000 2.69700000 ;
     RECT 7.73000000 2.47700000 7.95000000 2.69700000 ;
     RECT 8.85000000 2.47700000 9.07000000 2.69700000 ;
     RECT 9.97000000 2.47700000 10.19000000 2.69700000 ;
     RECT 11.09000000 2.47700000 11.31000000 2.69700000 ;
     RECT 12.21000000 2.47700000 12.43000000 2.69700000 ;
     RECT 13.33000000 2.47700000 13.55000000 2.69700000 ;
     RECT 14.45000000 2.47700000 14.67000000 2.69700000 ;
     RECT 15.57000000 2.47700000 15.79000000 2.69700000 ;
     RECT 16.69000000 2.47700000 16.91000000 2.69700000 ;
     RECT 17.81000000 2.47700000 18.03000000 2.69700000 ;
     RECT 18.93000000 2.47700000 19.15000000 2.69700000 ;
     RECT 1.01000000 2.88200000 1.23000000 3.10200000 ;
     RECT 2.13000000 2.88200000 2.35000000 3.10200000 ;
     RECT 3.25000000 2.88200000 3.47000000 3.10200000 ;
     RECT 4.37000000 2.88200000 4.59000000 3.10200000 ;
     RECT 5.49000000 2.88200000 5.71000000 3.10200000 ;
     RECT 6.61000000 2.88200000 6.83000000 3.10200000 ;
     RECT 7.73000000 2.88200000 7.95000000 3.10200000 ;
     RECT 8.85000000 2.88200000 9.07000000 3.10200000 ;
     RECT 9.97000000 2.88200000 10.19000000 3.10200000 ;
     RECT 11.09000000 2.88200000 11.31000000 3.10200000 ;
     RECT 12.21000000 2.88200000 12.43000000 3.10200000 ;
     RECT 13.33000000 2.88200000 13.55000000 3.10200000 ;
     RECT 14.45000000 2.88200000 14.67000000 3.10200000 ;
     RECT 15.57000000 2.88200000 15.79000000 3.10200000 ;
     RECT 16.69000000 2.88200000 16.91000000 3.10200000 ;
     RECT 17.81000000 2.88200000 18.03000000 3.10200000 ;
     RECT 18.93000000 2.88200000 19.15000000 3.10200000 ;

    LAYER pdiffc ;
     RECT 19.61500000 3.27200000 19.86500000 3.52200000 ;
     RECT 0.29500000 4.48700000 0.54500000 4.73700000 ;

    LAYER ndiffc ;
     RECT 0.29500000 0.30200000 0.54500000 0.55200000 ;
     RECT 4.91500000 0.30200000 5.16500000 0.55200000 ;
     RECT 9.39500000 0.30200000 9.64500000 0.55200000 ;
     RECT 13.87500000 0.30200000 14.12500000 0.55200000 ;
     RECT 18.35500000 0.30200000 18.60500000 0.55200000 ;
     RECT 2.67500000 0.57200000 2.92500000 0.82200000 ;
     RECT 7.15500000 0.57200000 7.40500000 0.82200000 ;
     RECT 11.63500000 0.57200000 11.88500000 0.82200000 ;
     RECT 16.11500000 0.57200000 16.36500000 0.82200000 ;
     RECT 19.61500000 1.92200000 19.86500000 2.17200000 ;

    LAYER met1 ;
     RECT 0.00000000 -0.24000000 20.16000000 0.24000000 ;
     RECT 0.21500000 0.24000000 0.62500000 0.63200000 ;
     RECT 4.83500000 0.24000000 5.24500000 0.63200000 ;
     RECT 9.31500000 0.24000000 9.72500000 0.63200000 ;
     RECT 13.79500000 0.24000000 14.20500000 0.63200000 ;
     RECT 18.27500000 0.24000000 18.68500000 0.63200000 ;
     RECT 2.59500000 0.49200000 3.00500000 0.90200000 ;
     RECT 7.07500000 0.49200000 7.48500000 0.90200000 ;
     RECT 11.55500000 0.49200000 11.96500000 0.90200000 ;
     RECT 16.03500000 0.49200000 16.44500000 0.90200000 ;
     RECT 19.53500000 1.84200000 19.94500000 2.25200000 ;
     RECT 0.93000000 2.39700000 1.31000000 2.77700000 ;
     RECT 2.05000000 2.39700000 2.43000000 2.77700000 ;
     RECT 3.17000000 2.39700000 3.55000000 2.77700000 ;
     RECT 4.29000000 2.39700000 4.67000000 2.77700000 ;
     RECT 5.41000000 2.39700000 5.79000000 2.77700000 ;
     RECT 6.53000000 2.39700000 6.91000000 2.77700000 ;
     RECT 7.65000000 2.39700000 8.03000000 2.77700000 ;
     RECT 8.77000000 2.39700000 9.15000000 2.77700000 ;
     RECT 9.89000000 2.39700000 10.27000000 2.77700000 ;
     RECT 11.01000000 2.39700000 11.39000000 2.77700000 ;
     RECT 12.13000000 2.39700000 12.51000000 2.77700000 ;
     RECT 13.25000000 2.39700000 13.63000000 2.77700000 ;
     RECT 14.37000000 2.39700000 14.75000000 2.77700000 ;
     RECT 15.49000000 2.39700000 15.87000000 2.77700000 ;
     RECT 16.61000000 2.39700000 16.99000000 2.77700000 ;
     RECT 17.73000000 2.39700000 18.11000000 2.77700000 ;
     RECT 18.85000000 2.39700000 19.23000000 2.77700000 ;
     RECT 0.93000000 2.80200000 1.31000000 3.18200000 ;
     RECT 2.05000000 2.80200000 2.43000000 3.18200000 ;
     RECT 3.17000000 2.80200000 3.55000000 3.18200000 ;
     RECT 4.29000000 2.80200000 4.67000000 3.18200000 ;
     RECT 5.41000000 2.80200000 5.79000000 3.18200000 ;
     RECT 6.53000000 2.80200000 6.91000000 3.18200000 ;
     RECT 7.65000000 2.80200000 8.03000000 3.18200000 ;
     RECT 8.77000000 2.80200000 9.15000000 3.18200000 ;
     RECT 9.89000000 2.80200000 10.27000000 3.18200000 ;
     RECT 11.01000000 2.80200000 11.39000000 3.18200000 ;
     RECT 12.13000000 2.80200000 12.51000000 3.18200000 ;
     RECT 13.25000000 2.80200000 13.63000000 3.18200000 ;
     RECT 14.37000000 2.80200000 14.75000000 3.18200000 ;
     RECT 15.49000000 2.80200000 15.87000000 3.18200000 ;
     RECT 16.61000000 2.80200000 16.99000000 3.18200000 ;
     RECT 17.73000000 2.80200000 18.11000000 3.18200000 ;
     RECT 18.85000000 2.80200000 19.23000000 3.18200000 ;
     RECT 19.53500000 3.19200000 19.94500000 3.60200000 ;
     RECT 0.21500000 4.40700000 0.62500000 4.80000000 ;
     RECT 0.00000000 4.80000000 20.16000000 5.28000000 ;

    LAYER via1 ;
     RECT 2.67000000 0.56700000 2.93000000 0.82700000 ;
     RECT 7.15000000 0.56700000 7.41000000 0.82700000 ;
     RECT 11.63000000 0.56700000 11.89000000 0.82700000 ;
     RECT 16.11000000 0.56700000 16.37000000 0.82700000 ;
     RECT 19.61000000 1.91700000 19.87000000 2.17700000 ;
     RECT 0.99000000 2.45700000 1.25000000 2.71700000 ;
     RECT 2.11000000 2.45700000 2.37000000 2.71700000 ;
     RECT 3.23000000 2.45700000 3.49000000 2.71700000 ;
     RECT 4.35000000 2.45700000 4.61000000 2.71700000 ;
     RECT 5.47000000 2.45700000 5.73000000 2.71700000 ;
     RECT 6.59000000 2.45700000 6.85000000 2.71700000 ;
     RECT 7.71000000 2.45700000 7.97000000 2.71700000 ;
     RECT 8.83000000 2.45700000 9.09000000 2.71700000 ;
     RECT 9.95000000 2.45700000 10.21000000 2.71700000 ;
     RECT 11.07000000 2.45700000 11.33000000 2.71700000 ;
     RECT 12.19000000 2.45700000 12.45000000 2.71700000 ;
     RECT 13.31000000 2.45700000 13.57000000 2.71700000 ;
     RECT 14.43000000 2.45700000 14.69000000 2.71700000 ;
     RECT 15.55000000 2.45700000 15.81000000 2.71700000 ;
     RECT 16.67000000 2.45700000 16.93000000 2.71700000 ;
     RECT 17.79000000 2.45700000 18.05000000 2.71700000 ;
     RECT 18.91000000 2.45700000 19.17000000 2.71700000 ;
     RECT 0.99000000 2.86200000 1.25000000 3.12200000 ;
     RECT 2.11000000 2.86200000 2.37000000 3.12200000 ;
     RECT 3.23000000 2.86200000 3.49000000 3.12200000 ;
     RECT 4.35000000 2.86200000 4.61000000 3.12200000 ;
     RECT 5.47000000 2.86200000 5.73000000 3.12200000 ;
     RECT 6.59000000 2.86200000 6.85000000 3.12200000 ;
     RECT 7.71000000 2.86200000 7.97000000 3.12200000 ;
     RECT 8.83000000 2.86200000 9.09000000 3.12200000 ;
     RECT 9.95000000 2.86200000 10.21000000 3.12200000 ;
     RECT 11.07000000 2.86200000 11.33000000 3.12200000 ;
     RECT 12.19000000 2.86200000 12.45000000 3.12200000 ;
     RECT 13.31000000 2.86200000 13.57000000 3.12200000 ;
     RECT 14.43000000 2.86200000 14.69000000 3.12200000 ;
     RECT 15.55000000 2.86200000 15.81000000 3.12200000 ;
     RECT 16.67000000 2.86200000 16.93000000 3.12200000 ;
     RECT 17.79000000 2.86200000 18.05000000 3.12200000 ;
     RECT 18.91000000 2.86200000 19.17000000 3.12200000 ;
     RECT 19.61000000 3.26700000 19.87000000 3.52700000 ;

    LAYER met2 ;
     RECT 0.89000000 2.35700000 1.35000000 3.22200000 ;
     RECT 2.01000000 2.35700000 2.47000000 3.22200000 ;
     RECT 3.13000000 2.35700000 3.59000000 3.22200000 ;
     RECT 4.25000000 2.35700000 4.71000000 3.22200000 ;
     RECT 5.37000000 2.35700000 5.83000000 3.22200000 ;
     RECT 6.49000000 2.35700000 6.95000000 3.22200000 ;
     RECT 7.61000000 2.35700000 8.07000000 3.22200000 ;
     RECT 8.73000000 2.35700000 9.19000000 3.22200000 ;
     RECT 9.85000000 2.35700000 10.31000000 3.22200000 ;
     RECT 10.97000000 2.35700000 11.43000000 3.22200000 ;
     RECT 12.09000000 2.35700000 12.55000000 3.22200000 ;
     RECT 13.21000000 2.35700000 13.67000000 3.22200000 ;
     RECT 14.33000000 2.35700000 14.79000000 3.22200000 ;
     RECT 15.45000000 2.35700000 15.91000000 3.22200000 ;
     RECT 16.57000000 2.35700000 17.03000000 3.22200000 ;
     RECT 17.69000000 2.35700000 18.15000000 3.22200000 ;
     RECT 2.57000000 0.46700000 3.03000000 0.55700000 ;
     RECT 7.05000000 0.46700000 7.51000000 0.55700000 ;
     RECT 11.53000000 0.46700000 11.99000000 0.55700000 ;
     RECT 16.01000000 0.46700000 16.47000000 0.55700000 ;
     RECT 2.57000000 0.55700000 19.18000000 0.83700000 ;
     RECT 2.57000000 0.83700000 3.03000000 0.92700000 ;
     RECT 7.05000000 0.83700000 7.51000000 0.92700000 ;
     RECT 11.53000000 0.83700000 11.99000000 0.92700000 ;
     RECT 16.01000000 0.83700000 16.47000000 0.92700000 ;
     RECT 18.90000000 0.83700000 19.18000000 2.35700000 ;
     RECT 18.81000000 2.35700000 19.27000000 3.22200000 ;
     RECT 19.51000000 1.81700000 19.97000000 2.27700000 ;
     RECT 19.60000000 2.27700000 19.88000000 3.16700000 ;
     RECT 19.51000000 3.16700000 19.97000000 3.62700000 ;

 END
END MUX8

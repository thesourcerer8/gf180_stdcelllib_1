VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO MUX8
  CLASS CORE ;
  FOREIGN MUX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 20.150 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 20.150 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 20.150 0.250 ;
    END
  END VGND
  PIN Z
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 19.500 3.150 19.950 3.650 ;
        RECT 19.600 2.300 19.900 3.150 ;
        RECT 19.500 1.800 19.950 2.300 ;
    END
  END Z
  PIN IN4
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 13.200 2.350 13.650 3.200 ;
    END
  END IN4
  PIN S0
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 3.150 2.350 3.600 3.200 ;
    END
  END S0
  PIN IN0
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 4.250 2.350 4.700 3.200 ;
    END
  END IN0
  PIN S5
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 15.450 2.350 15.900 3.200 ;
    END
  END S5
  PIN S7
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 2.350 2.450 3.200 ;
    END
  END S7
  PIN IN5
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 14.350 2.350 14.800 3.200 ;
    END
  END IN5
  PIN IN1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.750 2.350 9.200 3.200 ;
    END
  END IN1
  PIN S1
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 7.600 2.350 8.050 3.200 ;
    END
  END S1
  PIN S3
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 6.500 2.350 6.950 3.200 ;
    END
  END S3
  PIN S6
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 10.950 2.350 11.450 3.200 ;
    END
  END S6
  PIN S2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 16.550 2.350 17.050 3.200 ;
    END
  END S2
  PIN IN2
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 17.700 2.350 18.150 3.200 ;
    END
  END IN2
  PIN IN3
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 5.350 2.350 5.850 3.200 ;
    END
  END IN3
  PIN IN7
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.350 1.350 3.200 ;
    END
  END IN7
  PIN S4
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 12.100 2.350 12.550 3.200 ;
    END
  END S4
  PIN IN6
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 9.850 2.350 10.300 3.200 ;
    END
  END IN6
END MUX8
END LIBRARY


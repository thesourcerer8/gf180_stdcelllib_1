VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ASYNC3
  CLASS CORE ;
  FOREIGN ASYNC3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.950 BY 5.050 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 4.800 8.950 5.300 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0.000 -0.250 8.950 0.250 ;
    END
  END VGND
  PIN CN
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 1.450 2.050 1.900 2.150 ;
        RECT 7.600 2.050 8.050 2.150 ;
        RECT 1.450 1.750 8.050 2.050 ;
        RECT 1.450 1.700 1.900 1.750 ;
        RECT 7.600 1.700 8.050 1.750 ;
    END
  END CN
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 8.300 3.150 8.750 3.650 ;
        RECT 5.350 2.750 5.850 2.800 ;
        RECT 8.400 2.750 8.700 3.150 ;
        RECT 5.350 2.450 8.700 2.750 ;
        RECT 5.350 2.350 5.850 2.450 ;
        RECT 8.400 2.300 8.700 2.450 ;
        RECT 8.300 1.800 8.750 2.300 ;
    END
  END C
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 0.900 2.750 1.350 3.200 ;
        RECT 3.150 2.750 3.600 2.800 ;
        RECT 0.900 2.450 3.600 2.750 ;
        RECT 0.900 2.350 1.350 2.450 ;
        RECT 3.150 2.350 3.600 2.450 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal2 ;
        RECT 2.000 3.400 2.450 3.500 ;
        RECT 6.500 3.400 6.950 3.500 ;
        RECT 2.000 3.100 6.950 3.400 ;
        RECT 2.000 3.050 2.450 3.100 ;
        RECT 6.500 3.050 6.950 3.100 ;
    END
  END B
END ASYNC3
END LIBRARY

